ac test
R1 1 2 2
L1 2 3 1m
C1 3 0 3u
VS 1 0 AC=10V 90
.ac LOG 10000 1 100MHZ
.end