*netlist example 2
R1 1 0 5
G2 1 0 1 2 2
R3 1 2 6
R4 2 0 8
vin 1 0 5
.op
.dc vin 0.25 5.0 0.25
.end