diode test
VS 1 0 5V
D1 1 0 DMOD 1
.dc VS 0.25 5.0 0.25
.end