*tran rc
VS 1 0 PULSE 0.1 1V 2ns 3ns 4ns 5ns 20ns
R1 1 2 1
L1 2 3 1m
C1 3 0 1u
.tran 1ns 1us
.end
