*netlist example 1
R1 1 0 5
G2 1 0 1 2 2
R3 1 2 6
R4 2 0 8
Is 0 2 10
.op
.end