dc_sweep_test
vin 1 0 5
R1 1 0 1
.dc vin 0.25 5.0 0.25
.end
