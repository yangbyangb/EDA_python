tran test
C1 1 0 1uF
VS 1 0 PULSE 0 1V 2ns 3ns 4ns 5ns 20ns
.op
.tran 1ns 1us
.end
